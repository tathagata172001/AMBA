module 
int a;
endmodule
